module uart_top
(

input clk

);

endmodule
